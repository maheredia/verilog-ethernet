


module tcp_tx
#(

)
tcp_tx_inst
(
  input             clk              ,
  input             rst_n            ,
  //Control:
  input             syn_send         ,
  input             ack_send         ,
  input             fin_send         ,
  //Datapath: TODO
);

endmodule